//------------------------------------------------------------------------
// Input Conditioner
//    1) Synchronizes input to clock domain
//    2) Debounces input
//    3) Creates pulses at edge transitions
//------------------------------------------------------------------------

module inputconditioner
(
input 	    clk,            // Clock domain to synchronize input to
input	    noisysignal,    // (Potentially) noisy input signal
output wire conditioned,    // Conditioned output signal
output reg  positiveedge,   // 1 clk pulse at rising edge of conditioned
output reg  negativeedge    // 1 clk pulse at falling edge of conditioned
);
    debouncer deb(clk, noisysignal, conditioned);

    reg prevconditioned = 0;
    always @(posedge clk ) begin
        if(conditioned == 0 & prevconditioned == 1) begin
            positiveedge <= 1;
        end
        else begin
            negativeedge <= 0;
        end
    end
endmodule

// only changes the input signal after it is stable for a given waittime
module debouncer
(
input       clk,   // Clock domain to synchronize input to
input       sig,   // (Potentially) noisy input signal
output reg  out    // Debounced output signal
);

    parameter counterwidth = 3; // Counter size, in bits, >= log2(waittime)
    parameter waittime = 2;     // Debounce delay, in clock cycles

    reg[counterwidth-1:0] counter = 0;
    reg synchronizer0 = 0;
    reg synchronizer1 = 0;

    //0 0 0 0 1 0 1 1 1 1
    always @(posedge clk ) begin
        // Case 1: previous signal is same as current output
        if(out == synchronizer1)
            counter <= 0;
        else begin
            // Case 2: Counter reaches maximum limit
            if( counter == waittime) begin
                counter <= 0;
                out <= synchronizer1;
            end
            // Case 3: Counter has not reached max limit
            else
                counter <= counter+1;
        end
        synchronizer0 <= sig;
        synchronizer1 <= synchronizer0;
    end
endmodule
